`include "g2bnbit.v"
module tb;
	parameter N=10;
	reg [N-1:0]g;
	wire [N-1:0]b;
	g2bnbit dut(.b(b),.g(g));
	initial begin
		$display("%0d bit grey to binary code converter",N);
		$monitor("g=%b, b=%b",g,b);
		repeat(10) begin
			g = $random;
			#1;
		end
	end
endmodule
// 10 bit grey to binary code converter
//# g=0100100100, b=0111000111
//# g=1010000001, b=1100000001
//# g=1000001001, b=1111110001
//# g=1001100011, b=1110111101
//# g=1100001101, b=1000001001
//# g=0110001101, b=0100001001
//# g=0001100101, b=0001000110
//# g=1000010010, b=1111100011
//# g=1100000001, b=1000000001
//# g=0100001101, b=0111110110
//
//# 10 bit grey to binary code converter
//# g=0100100100, b=0111000111
//# g=1010000001, b=1100000001
//# g=1000001001, b=1111110001
//# g=1001100011, b=1110111101
//# g=1100001101, b=1000001001
//# g=0110001101, b=0100001001
//# g=0001100101, b=0001000110
//# g=1000010010, b=1111100011
//# g=1100000001, b=1000000001
//# g=0100001101, b=0111110110
