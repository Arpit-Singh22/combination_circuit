`include "encoder83.v"
module tb_encoder83;
	reg [7:0]i;
	wire [2:0]y;

	encoder83 dut(.i(i),.y(y));
	initial begin
		$monitor("i=%b, y=%b",i,y);
		i=8'b0000_0001;
		#1;
		i=8'b0000_0010;
		#1;
		i=8'b0000_0100;
		#1;
		i=8'b0000_1000;
		#1;
		i=8'b0001_0000;
		#1;
		i=8'b0001_0000;
		#1;
		i=8'b0010_0000;
		#1;
		i=8'b0100_0000;
		#1;
		i=8'b1000_0000;
		#1;
		i=8'b0010_0001;
		#1;	
	end
endmodule
//# i=00000001, y=000
//# i=00000010, y=001
//# i=00000100, y=010
//# i=00001000, y=011
//# i=00010000, y=100
//# i=00100000, y=101
//# i=01000000, y=110
//# i=10000000, y=111
//# i=00100001, y=zzz
